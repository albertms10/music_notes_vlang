module note

pub enum BaseNote {
	c = 0
	d = 2
	e = 4
	f = 5
	g = 7
	a = 9
	b = 11
}
